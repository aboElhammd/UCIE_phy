module SB_RX_HEADER_DECODER (
	input 				i_clk,
	input 				i_rst_n,
	input 				i_start_EN,
	input		[63:0]  i_header,
	output 	reg			o_tx_point_sweep_test_en,
	output 	reg	[1:0]  	o_tx_point_sweep_test,
	output 	reg	[3:0]	o_msg_no,
	output 	reg	[2:0]	o_msg_info,
	output 	reg			o_dec_header_valid
);


reg 	[1:0] 	test_type_reg;
wire 	[7:0] 	MsgCode;
wire 	[7:0] 	MsgSubCode;
wire 	[4:0]  	Opcode;
wire 	[15:0] 	MsgInfo;

assign Opcode 		= i_header [4:0];
assign MsgCode 		= i_header [21:14];
assign MsgSubCode 	= i_header [39:32];
assign MsgInfo 		= i_header [55:40];


//////////////////////////////////////////////////
/////// Point / Sweep Tests Enable And Test No.
//////////////////////////////////////////////////
always @(posedge i_clk or negedge i_rst_n) begin
	if(~i_rst_n) begin
		o_tx_point_sweep_test_en	<= 0;
		o_tx_point_sweep_test 		<= 0;
	end 
	else if (i_start_EN) begin
		if (MsgCode [7:4] == 4'h8) begin
			o_tx_point_sweep_test_en <= 1;
			case (MsgSubCode)
				8'h01: o_tx_point_sweep_test <= 00;
				8'h05: o_tx_point_sweep_test <= 01;
				8'h07: o_tx_point_sweep_test <= 10;
				8'h0A: o_tx_point_sweep_test <= 11;
			endcase

		end
		else begin
			o_tx_point_sweep_test_en <= 0;
		end
	end
	/*else begin
		o_tx_point_sweep_test_en <= 0;
	end*/
end


//////////////////////////////////////////////////
/////// MsgNo and MsgInfo
//////////////////////////////////////////////////
always @(posedge i_clk or negedge i_rst_n) begin
	if(~i_rst_n) begin
		o_msg_no 				<= 0;
		o_msg_info 				<= 0;
	end 
	else if (i_start_EN) begin
		if (MsgCode [7:4] == 4'h8) begin
			case (MsgSubCode)
				8'h01, 8'h05, 8'h07, 8'h0A://------------------------------------------------------------------------------
				  	begin
				  		case (MsgCode [3:0])
				  			4'h5://------------------------------------------------------------------------------
				  				begin
				  					o_msg_no  	<= 1;
				  					//o_msg_info 	<= ??; //******************
 				  				end
				  			//------------------------------------------------------------------------------
				  			4'hA://------------------------------------------------------------------------------
				  				begin
				  					o_msg_no  	<= 2;
				  					o_msg_info 	<= 0; //******************
 				  				end
				  			//------------------------------------------------------------------------------
				  		endcase
				  	end
				//------------------------------------------------------------------------------
			
				8'h02://------------------------------------------------------------------------------
				  	begin
				  		o_msg_info 	<= 0;
				  		case (MsgCode [3:0])
				  			4'h5://------------------------------------------------------------------------------
				  				begin
				  					o_msg_no  	<= 3;
 				  				end
				  			//------------------------------------------------------------------------------
				  			4'hA://------------------------------------------------------------------------------
				  				begin
				  					o_msg_no  	<= 4;
 				  				end
				  			//------------------------------------------------------------------------------
				  		endcase
				  	end
				//------------------------------------------------------------------------------
			
				8'h03, 8'h0B://------------------------------------------------------------------------------
				  	begin
				  		case (MsgCode [3:0])
				  			4'h5://------------------------------------------------------------------------------
				  				begin
				  					o_msg_no  	<= 5;
				  					o_msg_info 	<= 0;
 				  				end
				  			//------------------------------------------------------------------------------
				  			4'hA://------------------------------------------------------------------------------
				  				begin
				  					o_msg_no  	<= 6;
				  					//o_msg_info 	<= ??; //******************
 				  				end
				  			//------------------------------------------------------------------------------
				  		endcase
				  	end
				//------------------------------------------------------------------------------

				8'h04, 8'h09, 8'h0D://------------------------------------------------------------------------------
				  	begin
				  		o_msg_info 	<= 0;
				  		case (MsgCode [3:0])
				  			4'h5://------------------------------------------------------------------------------
				  				begin
				  					o_msg_no  	<= 7;
 				  				end
				  			//------------------------------------------------------------------------------
				  			4'hA://------------------------------------------------------------------------------
				  				begin
				  					o_msg_no  	<= 8;
 				  				end
				  			//------------------------------------------------------------------------------
				  		endcase
				  	end
				//------------------------------------------------------------------------------

				8'h06, 8'h08://------------------------------------------------------------------------------
				  	begin
				  		o_msg_info 	<= 0;
				  		case (MsgCode [3:0])
				  			4'h5://------------------------------------------------------------------------------
				  				begin
				  					o_msg_no  	<= 5;
 				  				end
				  			//------------------------------------------------------------------------------
				  			4'hA://------------------------------------------------------------------------------
				  				begin
				  					o_msg_no  	<= 6;
 				  				end
				  			//------------------------------------------------------------------------------
				  		endcase
				  	end
				//------------------------------------------------------------------------------

				8'h0C://------------------------------------------------------------------------------
					begin
						o_msg_no 	<= 9;
						o_msg_info 	<= 0;
					end
				//------------------------------------------------------------------------------			
			endcase
		end
		
		else if (MsgCode [7:4] == 4'h9) begin
			case (MsgSubCode)
				8'h00://------------------------------------------------------------------------------
					begin
						o_msg_no 	<= 3;
						o_msg_info 	<= 0;
					end
				//------------------------------------------------------------------------------			
			
				8'h01://------------------------------------------------------------------------------
					begin
						o_msg_info 	<= 0;
						case (MsgCode [3:0])
							4'h5://------------------------------------------------------------------------------
								begin
									o_msg_no 	<= 1;
								end
							//------------------------------------------------------------------------------

							4'hA://------------------------------------------------------------------------------
								begin
									o_msg_no 	<= 2;
								end
							//------------------------------------------------------------------------------	
						endcase
					end
				//------------------------------------------------------------------------------

			endcase
		end
		
		else if (MsgCode [7:4] == 4'hA) begin
			case (MsgSubCode)
				8'h00,8'h02,8'h03,8'h09,8'h0D,8'h11://------------------------------------------------------------------------------1 -	2	-	msginfo = 0
					begin
						o_msg_info 	<= 0;
						case (MsgCode [3:0])
							4'h5://------------------------------------------------------------------------------
								begin
									o_msg_no 	<= 1;
								end
							//------------------------------------------------------------------------------

							4'hA://------------------------------------------------------------------------------
								begin
									o_msg_no 	<= 2;
								end
							//------------------------------------------------------------------------------	
						endcase
					end
				//------------------------------------------------------------------------------

				8'h04,8'h0A://------------------------------------------------------------------------------3 -	4	-	msginfo != 0
					begin
						case (MsgCode [3:0])
							4'h5://------------------------------------------------------------------------------
								begin
									o_msg_no 	<= 3;
									o_msg_info 	<= 0;
								end
							//------------------------------------------------------------------------------

							4'hA://------------------------------------------------------------------------------
								begin
									o_msg_no 	<= 4;
									o_msg_info 	<= MsgInfo[2:0];
								end
							//------------------------------------------------------------------------------	
						endcase
					end
				//------------------------------------------------------------------------------

				8'h08,8'h0C,8'h0F://------------------------------------------------------------------------------5 -	6	-	msginfo = 0
					begin
						o_msg_info 	<= 0;
						case (MsgCode [3:0])
							4'h5://------------------------------------------------------------------------------
								begin
									o_msg_no 	<= 5;
								end
							//------------------------------------------------------------------------------

							4'hA://------------------------------------------------------------------------------
								begin
									o_msg_no 	<= 6;
								end
							//------------------------------------------------------------------------------	
						endcase
					end
				//------------------------------------------------------------------------------

				

				8'h0E,8'h13://------------------------------------------------------------------------------3 -	4	-	msginfo = 0
					begin
						o_msg_info 	<= 0;
						case (MsgCode [3:0])
							4'h5://------------------------------------------------------------------------------
								begin
									o_msg_no 	<= 3;
								end
							//------------------------------------------------------------------------------

							4'hA://------------------------------------------------------------------------------
								begin
									o_msg_no 	<= 4;
								end
							//------------------------------------------------------------------------------	
						endcase
					end
				//------------------------------------------------------------------------------

				8'h10://------------------------------------------------------------------------------7 -	8	-	msginfo = 0
					begin
						o_msg_info 	<= 0;
						case (MsgCode [3:0])
							4'h5://------------------------------------------------------------------------------
								begin
									o_msg_no 	<= 7;
								end
							//------------------------------------------------------------------------------

							4'hA://------------------------------------------------------------------------------
								begin
									o_msg_no 	<= 8;
								end
							//------------------------------------------------------------------------------	
						endcase
					end
				//------------------------------------------------------------------------------

				8'h14://------------------------------------------------------------------------------5 -	6	-	msginfo != 0
					begin
						case (MsgCode [3:0])
							4'h5://------------------------------------------------------------------------------
								begin
									o_msg_no 	<= 5;
									o_msg_info 	<= MsgInfo[2:0];
								end
							//------------------------------------------------------------------------------

							4'hA://------------------------------------------------------------------------------
								begin
									o_msg_no 	<= 6;
									o_msg_info 	<= 0;
								end
							//------------------------------------------------------------------------------	
						endcase
					end
				//-----------------------------------------------------------------------------
			endcase
		end

		else if (MsgCode [7:4] == 4'hB) begin
			case (MsgSubCode)
				8'h00,8'h02,8'h04,8'h05,8'h06,8'h08,8'h0A,8'h0C,8'h0E,8'h11,8'h13,8'h15,8'h1B://------------------------------------------------------------------------------1 -	2	-	msginfo = 0
					begin
						o_msg_info 	<= 0;
						case (MsgCode [3:0])
							4'h5://------------------------------------------------------------------------------
								begin
									o_msg_no 	<= 1;
								end
							//------------------------------------------------------------------------------

							4'hA://------------------------------------------------------------------------------
								begin
									o_msg_no 	<= 2;
								end
							//------------------------------------------------------------------------------	
						endcase
					end
				//------------------------------------------------------------------------------

				8'h01,8'h03,8'h07,8'h09,8'h0B,8'h0D,8'h10,8'h12,8'h14,8'h16,8'h1C://------------------------------------------------------------------------------3 -	4	-	msginfo = 0
					begin
						o_msg_info 	<= 0;
						case (MsgCode [3:0])
							4'h5://------------------------------------------------------------------------------
								begin
									o_msg_no 	<= 3;
								end
							//------------------------------------------------------------------------------

							4'hA://------------------------------------------------------------------------------
								begin
									o_msg_no 	<= 4;
								end
							//------------------------------------------------------------------------------	
						endcase
					end
				//------------------------------------------------------------------------------			

				8'h17,8'h1D://------------------------------------------------------------------------------5 -	6	-	msginfo = 0
					begin
						o_msg_info 	<= 0;
						case (MsgCode [3:0])
							4'h5://------------------------------------------------------------------------------
								begin
									o_msg_no 	<= 5;
								end
							//------------------------------------------------------------------------------

							4'hA://------------------------------------------------------------------------------
								begin
									o_msg_no 	<= 6;
								end
							//------------------------------------------------------------------------------	
						endcase
					end
				//------------------------------------------------------------------------------

				8'h18://------------------------------------------------------------------------------7 -	8	-	msginfo = 0
					begin
						o_msg_info 	<= 0;
						case (MsgCode [3:0])
							4'h5://------------------------------------------------------------------------------
								begin
									o_msg_no 	<= 7;
								end
							//------------------------------------------------------------------------------

							4'hA://------------------------------------------------------------------------------
								begin
									o_msg_no 	<= 8;
								end
							//------------------------------------------------------------------------------	
						endcase
					end
				//------------------------------------------------------------------------------

				8'h1E://------------------------------------------------------------------------------7 -	8	-	msginfo != 0
					begin
						case (MsgCode [3:0])
							4'h5://------------------------------------------------------------------------------
								begin
									o_msg_no 	<= 7;
									o_msg_info 	<= MsgInfo[2:0];
								end
							//------------------------------------------------------------------------------

							4'hA://------------------------------------------------------------------------------
								begin
									o_msg_no 	<= 8;
									o_msg_info 	<= 0;
								end
							//------------------------------------------------------------------------------	
						endcase
					end
				//------------------------------------------------------------------------------

				8'h19://------------------------------------------------------------------------------7 -	8	-	msginfo = 0
					begin
						o_msg_info 	<= 0;
						case (MsgCode [3:0])
							4'h5://------------------------------------------------------------------------------
								begin
									o_msg_no 	<= 9;
								end
							//------------------------------------------------------------------------------

							4'hA://------------------------------------------------------------------------------
								begin
									o_msg_no 	<= 10;
								end
							//------------------------------------------------------------------------------	
						endcase
					end
				//------------------------------------------------------------------------------

				8'h1F://------------------------------------------------------------------------------7 -	8	-	msginfo = 0
					begin
						o_msg_info 	<= 0;
						case (MsgCode [3:0])
							4'h5://------------------------------------------------------------------------------
								begin
									o_msg_no 	<= 11;
								end
							//------------------------------------------------------------------------------

							4'hA://------------------------------------------------------------------------------
								begin
									o_msg_no 	<= 12;
								end
							//------------------------------------------------------------------------------	
						endcase
					end
				//------------------------------------------------------------------------------



			endcase
		end

		else if (MsgCode [7:4] == 4'hC) begin
			case (MsgSubCode)
				8'h01://------------------------------------------------------------------------------1 -	2	-	msginfo = 0
					begin
						o_msg_info 	<= MsgInfo[2:0];
						case (MsgCode [3:0])
							4'h5://------------------------------------------------------------------------------
								begin
									o_msg_no 	<= 1;
								end
							//------------------------------------------------------------------------------

							4'hA://------------------------------------------------------------------------------
								begin
									o_msg_no 	<= 2;
								end
							//------------------------------------------------------------------------------	
						endcase
					end
				//------------------------------------------------------------------------------

			endcase
		end

		else if (MsgCode [7:4] == 4'hE) begin
			case (MsgSubCode)
				8'h00://------------------------------------------------------------------------------1 -	2	-	msginfo = 0
					begin
						o_msg_info 	<= 0;
						case (MsgCode [3:0])
							4'h5://------------------------------------------------------------------------------
								begin
									o_msg_no 	<= 15;
								end
							//------------------------------------------------------------------------------

							4'hA://------------------------------------------------------------------------------
								begin
									o_msg_no 	<= 14;
								end
							//------------------------------------------------------------------------------	
						endcase
					end
				//------------------------------------------------------------------------------

			endcase
		end

	end
end

//////////////////////////////////////////////////
/////// Output Valid
//////////////////////////////////////////////////
always @(posedge i_clk or negedge i_rst_n) begin
	if(~i_rst_n) begin
		o_dec_header_valid <= 0;
	end 
	else if (i_start_EN) begin
		o_dec_header_valid <= 1;
	end
	else if (o_dec_header_valid) begin
		o_dec_header_valid <= 0;
	end
end




endmodule : SB_RX_HEADER_DECODER


//////////////////////////////////////////////////
/////// Opcode Dencoding (Packet With/Without Data)
//////////////////////////////////////////////////
/*always @(posedge i_clk or negedge i_rst_n) begin
	if(~i_rst_n) begin
		o_packet_with_data <= 0;
	end 
	else if (i_start_EN) begin
		if (Opcode == 5'b11011) begin
			o_packet_with_data <= 1;
		end
		else begin
			o_packet_with_data <= 0;
		end
	end
	else if (o_packet_with_data) begin
		o_packet_with_data <= 0;
	end
end*/