module RX_TRAINERROR_HS #(
    parameter SB_MSG_WIDTH = 4
) (
    input                                        i_clk,
    input                                        i_rst_n, 
    input                                        i_trainerror_en,           // eli gyaly mn module el LTSM 34an abd2 asasn di el enable bta3t this module
	input 										 i_rx_msg_valid,
	input   									 i_falling_edge_busy,	    // gayly mn elSB 34an y2olii enu khalas ba3t el data bta3te fa anzl el valid
   	input   									 i_SB_Busy,		 		    // gayly mn elSB 34an y2olii enu khalas ba3t el data bta3te fa anzl el valid
	input 										 i_partner_req_trainerror,
    input                                        i_tx_valid,
    input       [SB_MSG_WIDTH-1:0]               i_decoded_SB_msg,          // gyaly mn el SB b3d my3ml decode ll msg eli gyalo mn el partner w yb3tli el crossponding format liha 
    output reg  [SB_MSG_WIDTH-1:0]               o_encoded_SB_msg_rx,       // sent to SB 34an 22olo haystkhdm anhy encoding
    output reg                                   o_trainerror_end_rx,       // sent to LTSM 34an ykhush el TRAINERROR w 22olo eni khalst
    output reg                                   o_valid_rx                 // sent to Wrapper 34an 22olo eni 3ndi data valid 3ayz ab3tha
);

/////////////////////////////////////////
//////////// Internal signals ///////////
/////////////////////////////////////////

reg [2:0] CS, NS; // Current State, Next State	

// dool el conditions eli batl3 el outputs based 3alehum
wire send_trainerror_entry_resp, send_trainerror_end;
reg save_resp_state;
reg save_rx_valid; // register used to detect the falling edge of the vaild to be used as a condition for transitions in next state logic

/////////////////////////////////////////
//////////// Machine STATES /////////////
/////////////////////////////////////////

localparam [2:0] IDLE     					    = 0;
localparam [2:0] WAIT_FOR_TRAINERROR_REQ        = 1;
localparam [2:0] SEND_TRAINERROR_RESP		    = 2;
localparam [2:0] TEST_FINISHED    				= 3;

/////////////////////////////////////////
///////////// SB messages ///////////////
/////////////////////////////////////////

localparam TRAINERROR_entry_req_msg 	= 15;
localparam TRAINERROR_entry_resp_msg	= 14;

/////////////////////////////////////////
////////// Assign statements ////////////
/////////////////////////////////////////

assign send_trainerror_entry_resp  = (CS == WAIT_FOR_TRAINERROR_REQ && NS == SEND_TRAINERROR_RESP); 
assign send_trainerror_end	       = (CS == SEND_TRAINERROR_RESP && NS == TEST_FINISHED );
wire   falling_edge_valid 		   = (save_rx_valid != o_valid_rx) && !o_valid_rx;

/////////////////////////////////
//////// State Memory ///////////
/////////////////////////////////

always @ (posedge i_clk or negedge i_rst_n) begin
    if (!i_rst_n) begin
        CS <= IDLE;
    end
    else begin
        CS <= NS;
    end
end

/////////////////////////////////
/////// Next State Logic ////////
/////////////////////////////////

always @ (*) begin
	case (CS) 
/*-----------------------------------------------------------------------------
* IDLE
*-----------------------------------------------------------------------------*/
		IDLE: begin
			NS = (i_trainerror_en)? WAIT_FOR_TRAINERROR_REQ   : IDLE;
		end
/*-----------------------------------------------------------------------------
* WAIT_FOR_TRAINERROR_REQ    
*-----------------------------------------------------------------------------*/
        WAIT_FOR_TRAINERROR_REQ  : begin 
            if (i_trainerror_en) begin
				if ((i_decoded_SB_msg == TRAINERROR_entry_req_msg && i_rx_msg_valid) || i_partner_req_trainerror) begin 
					NS = SEND_TRAINERROR_RESP;
				end 
				else begin
					NS = WAIT_FOR_TRAINERROR_REQ;
				end
            end else begin
                NS = IDLE;
            end
        end
/*-----------------------------------------------------------------------------
* SEND_TRAINERROR_RESP
*-----------------------------------------------------------------------------*/
		SEND_TRAINERROR_RESP: begin
            if (i_trainerror_en) begin
				if (falling_edge_valid) begin // m3anaha en el SB khalas khd el data mn 3al bus 
					NS = TEST_FINISHED;
				end 
				else begin
					NS = SEND_TRAINERROR_RESP;
				end
            end else begin
                NS = IDLE;
            end
		end
/*-----------------------------------------------------------------------------
* TEST_FINISHED 
*-----------------------------------------------------------------------------*/
		TEST_FINISHED   : begin
			if (!i_trainerror_en) begin
				NS = IDLE;
			end else begin
				NS = TEST_FINISHED;
			end
		end
		default: NS = IDLE;
    endcase
end

/////////////////////////////////
///////// Output Logic //////////
/////////////////////////////////

always @ (posedge i_clk or negedge i_rst_n) begin
    if (!i_rst_n) begin
        o_trainerror_end_rx <= 0;
        o_encoded_SB_msg_rx <= 0;
    end
    else begin
        if (CS == IDLE) begin
            o_trainerror_end_rx <= 0;
            o_encoded_SB_msg_rx <= 0;
        end
        
        if (send_trainerror_entry_resp) begin
            o_encoded_SB_msg_rx <= TRAINERROR_entry_resp_msg;
        end
        
        if (send_trainerror_end) begin
            o_trainerror_end_rx <= 1;
        end
    end
end

/////////////////////////////////
////////// Valid Logic //////////
/////////////////////////////////
always @(posedge i_clk or negedge i_rst_n ) begin
	if (!i_rst_n) begin
		o_valid_rx <= 0;
		save_rx_valid <= 0;
	end else begin
		save_rx_valid <= o_valid_rx;
		if (i_falling_edge_busy) begin 
			o_valid_rx <= 0;
		end
		else if ((send_trainerror_entry_resp && !i_SB_Busy) || (save_resp_state && !i_tx_valid)) begin  
			o_valid_rx <= 1;
		end
	end
end

always @ (posedge i_clk or negedge i_rst_n) begin
	if (!i_rst_n) begin
		save_resp_state <= 0;
	end else begin
		if (send_trainerror_entry_resp && i_tx_valid) begin
			save_resp_state <= 1; 
			// el flag dh ana 3amlo 34an lw el tx byb3t fa bltaly ana mynf34 arf3 el valid bta3 el rx bas fi nafs el w2t me7tag a save eni kunt me7tag arf3 elvalid
			// mn gher el flag dh el condition eli kan bykhlene arf3 elvalid eli hwa dh lw7do (send_done_rsp && !i_SB_Busy) kan 1 clock cycle w bydee3 fa bltaly 
			// mkunt4 ba3rf arf3 elvalid lakn dlwi2ty ana ba save eni elmafrood arf3 el valid b3d ma el tx ykhls mn khelal el flag dh
		end else if (o_valid_rx) begin
			save_resp_state <= 0;
		end
	end 
end 

endmodule